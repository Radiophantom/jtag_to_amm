
package amm_regs_pkg;

  parameter logic [15:0] REGS_RO_MASK [32] = '{
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF,
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF,
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF,
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF,
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF,
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF,
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF,
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF
  };

  parameter logic [15:0] REGS_INIT [32] = '{
    16'hAAAA,
    16'hBBBB,
    16'hCCCC,
    16'hDDDD,
    16'hAAAA,
    16'hBBBB,
    16'hCCCC,
    16'hDDDD,
    16'hAAAA,
    16'hBBBB,
    16'hCCCC,
    16'hDDDD,
    16'hAAAA,
    16'hBBBB,
    16'hCCCC,
    16'hDDDD,
    16'hAAAA,
    16'hBBBB,
    16'hCCCC,
    16'hDDDD,
    16'hAAAA,
    16'hBBBB,
    16'hCCCC,
    16'hDDDD,
    16'hAAAA,
    16'hBBBB,
    16'hCCCC,
    16'hDDDD,
    16'hAAAA,
    16'hBBBB,
    16'hCCCC,
    16'hDDDD
  };

endpackage

