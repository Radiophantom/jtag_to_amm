
package amm_regs_pkg;

  parameter bit [0:31][15:0] regs_ro_mask = {
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF,
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF,
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF,
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF,
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF,
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF,
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF,
    16'h0000,
    16'h00FF,
    16'hFF00,
    16'hFFFF
  };

  parameter bit [0:31][15:0] regs_init = {
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD,
    16'hABCD
  };

endpackage

